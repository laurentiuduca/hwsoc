// laur
`define SIM_MODE
`define TN_DRAM_REFRESH // for tang nano
`define SIM_TNSRAM // tang nano not only sim ram

`define FREQ 27_000_000
`define MEM_SIZE (8*1024*1024)
`define BBL_SIZE (8*1024*1024)

`define CACHE_SIZE (32*1024)

`define XLEN    32
`define LATENCY 0
